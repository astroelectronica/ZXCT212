.title KiCad schematic
.include "C:/AE/ZXCT212/CEU4J2X7R2A103K125AE_s.mod"
.include "C:/AE/ZXCT212/ZXCT212.LIB"
I1 /IN- 0 DC {ILOAD} 
XU2 /OUT 0 CEU4J2X7R2A103K125AE_s
R2 /CNV /OUT {ROUT}
R1 /IN- /VIN {RSNS}
XU1 /VREF 0 /VSUPPLY /VIN /IN- /CNV ZXCT212
V2 /VREF 0 DC {VREF} 
V1 /VIN 0 DC {VIN} 
V3 /VSUPPLY 0 DC {VSUPPLY} 
.end
